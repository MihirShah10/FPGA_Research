module jpeg ( 
input			clk ,			// line#=./dct.h:23
input			rst ,			// line#=./dct.h:24
input	[11:0]	jpeg_in_a00 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a01 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a02 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a03 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a04 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a05 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a06 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a07 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a08 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a09 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a10 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a11 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a12 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a13 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a14 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a15 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a16 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a17 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a18 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a19 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a20 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a21 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a22 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a23 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a24 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a25 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a26 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a27 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a28 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a29 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a30 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a31 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a32 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a33 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a34 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a35 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a36 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a37 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a38 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a39 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a40 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a41 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a42 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a43 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a44 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a45 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a46 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a47 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a48 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a49 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a50 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a51 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a52 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a53 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a54 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a55 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a56 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a57 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a58 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a59 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a60 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a61 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a62 ,	// line#=./dct.h:27
input	[11:0]	jpeg_in_a63 ,	// line#=./dct.h:27
output	[11:0]	jpeg_out_a00 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a01 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a02 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a03 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a04 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a05 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a06 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a07 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a08 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a09 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a10 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a11 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a12 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a13 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a14 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a15 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a16 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a17 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a18 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a19 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a20 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a21 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a22 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a23 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a24 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a25 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a26 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a27 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a28 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a29 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a30 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a31 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a32 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a33 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a34 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a35 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a36 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a37 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a38 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a39 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a40 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a41 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a42 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a43 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a44 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a45 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a46 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a47 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a48 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a49 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a50 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a51 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a52 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a53 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a54 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a55 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a56 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a57 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a58 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a59 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a60 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a61 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a62 ,	// line#=./dct.h:30
output	[11:0]	jpeg_out_a63 ,	// line#=./dct.h:30
output		    valid			// line#=./dct.h:31
);

endmodule